library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_Contador is
end tb_Contador;

architecture Behavioral of tb_Contador is

    -- Component Declaration for the Unit Under Test (UUT)
    component Contador is
        port (
            Clock   : in  std_logic;
            Reset   : in  std_logic;
            Control : in  std_logic;
            Start   : in  std_logic_vector(3 downto 0);
            Enable  : in  std_logic;
            Count   : out std_logic_vector(3 downto 0)
        );
    end component;

    -- Signals to connect to UUT
    signal Clock   : std_logic := '0';
    signal Reset   : std_logic := '0';
    signal Control : std_logic := '0';
    signal Start   : std_logic_vector(3 downto 0) := "0000";
    signal Enable  : std_logic := '0';
    signal Count   : std_logic_vector(3 downto 0);

    -- Clock period definition
    constant Clock_period : time := 10 ns;

begin

    -- Instantiate the Unit Under Test (UUT)
    uut: Contador
        port map (
            Clock   => Clock,
            Reset   => Reset,
            Control => Control,
            Start   => Start,
            Enable  => Enable,
            Count   => Count
        );

    -- Clock generation process
    Clock_process :process
    begin
        Clock <= '0';
        wait for Clock_period/2;
        Clock <= '1';
        wait for Clock_period/2;
    end process;

    -- Stimulus process
    stim_proc: process
    begin        
        -- hold reset state for 20 ns.
        wait for 20 ns;  
        Reset <= '1';
        wait for 20 ns;
        Reset <= '0';

        -- Test case 1: Enable and increment
        Start <= "0000";
        Control <= '1';
        Enable <= '1';
        wait for 20 ns;
        
        -- Test case 2: Disable and hold
        Enable <= '0';
        wait for 20 ns;

        -- Test case 3: Decrement
        Enable <= '1';
        Control <= '0';
        wait for 40 ns;
        
        -- Test case 4: Reset and start from a non-zero value
		  wait for 20 ns;
        Start <= "0100";
		  Reset <= '1';
		  wait for 20 ns;
        Reset <= '0';
        Control <= '1';
        wait for 100 ns;

        -- Stop simulation
        wait;
    end process;

end Behavioral;
